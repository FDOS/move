# Hjälpmeddelanden

0.0:Move
0.1:Flytter en fil/katalog till en annan plats.
0.2:(C) 1997-2002 by Joe Cosentino
0.3:(C) 2003-2004 by Imre Leber
0.4:Syntax: MOVE
0.5:källa1[, källa2[,...]] destination
0.6: källa       Namnet på filen eller katalogen du vill flytta (byta namn på)
0.7: destination Vart du vill flytta filen/filerna
0.8:          Undertrycker förfrågan om du vill skriva över
0.9:             en existerande destinations fil.
0.10:         Ser till att förfrågan sker om överskrivning av
0.11:             existerande destinationsfil.
0.12:          Verifierar varje file då den skrivs till destinationsfilen
0.13:             för att säkerställa att destinations filerna är identiska med
0.14:             källfilerna
0.15:Not:
0.16:Du kan flytta kataloger med detta verktyg

# Diverse meddelanden

1.0:finns ej!
1.1:finns redan!
1.2:Skriv över fil
1.3:Problem vid förflyttning av katalog
1.4:Problem vid förflyttning av fil
1.5:Ogiltig parameter
1.6:Ogiltig enhetsspecifikation för källa
1.7:Ogiltig destinationsfil
1.8: finns inte som en katalog. Skapa den?
1.9:Ogiltig källfil
1.10:Kan inte skapa katalog
1.11:Fil kan inte kopieras ovanpå sig själv
1.12:Kan inte flytta en fil till en katalog
1.13:Fil finns redan
1.14:Fil kan inte kopieras ovanpå sig själv
1.15:Åtkomst nekad
1.16:Otillräckligt diskutrymme i destinationssökväg
1.17:Otillräckligt diskutrymme
1.18:Nödvändig parameter saknas
1.19:Ogiltig källspecifikation
1.20:Källsökväg finns inte
1.21:Källsökväg för lång\n
1.22:Destinationssökväg för lång\n
1.23:Ogiltig enhetsspecifikation för destination\n
1.24:Destinationssökväg för lång\n
1.25:Kan inte öppna källfil
1.26:Kan inte skapa destinationsfil
1.27:Skrivfel vid destinationsfil
1.28:Kan inte skapa katalog
1.29:Otillräckligt diskutrymme i destinationssökväg

# J/N/Alla/Inga; Enkla meddelanden

2.0:J
2.1:N
2.2:Alla
2.3:Inga
2.4:ok
